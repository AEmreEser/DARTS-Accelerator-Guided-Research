`timescale 1ns/1ps
module PE_matrix_simple_tb;
   localparam int FILT_SIZE  = 3;
   localparam int PSUM_WIDTH = 36;

   logic  clk = 0;
   logic  rst = 1;

   logic  start;
   logic  done;
   
   logic signed [5:0] counter;

   logic signed [15:0] Filt [2:0][2:0];
   logic signed [15:0] Img  [27:0][27:0];
   logic [PSUM_WIDTH-1:0] output_psum       [25:0][25:0];
   logic [PSUM_WIDTH-1:0] output_psum_golden[25:0][25:0] = '{
    { 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000 },
    { 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000 },
    { 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000 },
    { 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000 },
    { 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000 },
    { 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000 },
    { 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000 },
    { 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000 },
    { 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000 },
    { 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000 },
    { 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000 },
    { 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000 },
    { 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000 },
    { 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000 },
    { 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000 },
    { 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000 },
    { 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000 },
    { 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000 },
    { 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000 },
    { 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000 },
    { 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000 },
    { 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000 },
    { 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000 },
    { 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000 },
    { 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000 },
    { 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000, 36'h000120000 }
};

   always #5ns clk = ~clk;

   PE_matrix #(.PSUM_WIDTH(PSUM_WIDTH)) pe_array_dut
   (
      .clk(clk),
      .rst(rst),
      .start(start),
      .rstAccumulation(1'b0),
      .Filt(Filt),
      .Img(Img),
      .counter(counter),
      .done(done),
      .output_psum(output_psum)
   );

   initial begin
      /* ---- stimuli ---- */
      

Filt = '{
    { 16'h0200, 16'h0200, 16'h0200 },
    { 16'h0200, 16'h0200, 16'h0200 },
    { 16'h0200, 16'h0200, 16'h0200 }
};

Img = '{
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 },
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 },
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 },
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 },
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 },
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 },
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 },
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 },
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 },
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 },
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 },
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 },
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 },
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 },
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 },
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 },
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 },
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 },
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 },
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 },
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 },
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 },
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 },
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 },
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 },
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 },
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 },
    { 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100 }
};

      /* reset sequence */
      rst   = 1'b1;
      start = 1'b0;
      repeat (2) @(negedge clk);
      rst   = 1'b0;

      /* single-cycle start pulse */
      @(negedge clk) start = 1'b1;
      @(negedge clk) start = 1'b0;

      if (done !== 1'b1) begin
         $display("Test failed: done signal not asserted as expected.");
         $finish;
      end
      #20000;

      $finish;
   end
endmodule
